module top_module( 
    input a, 
    input b, 
    output out );
    and (out,b,a);

endmodule