module top_module( input in, output out );
wire a;
    assign a = in;
    assign out = a;
endmodule